Complementaire Darlington met emitter degeneratie
*
*  PUSH-PULL TRANSISTOR OUTPUT STAGE
Q1 2 1 0 QNPN
Q2 0 2 3 QPNP
*
* DEVICE MODELS
.model QNPN	NPN(BF=50)
.model QPNP	PNP(BF=50)
* klasseF
Q_Q1         2 1 0 Q2
L_L1         0 3   1uH  
C_C1         0 3   10n  
R_R1         0 3   100  
V_V3         4 0   10V
V_V5         1 0   sin(0.4 0.8 1591500) DC=0.4
C_C3         5 3   10n  
L_L3         6 3   0.111uH
R_R3         6 5   0.001 
L_L2         2 4   2mH  
C_C2         2 5   1000n  
.model Q2  NPN(Is=14.34f BF=200 Rb=100 )

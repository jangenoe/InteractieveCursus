* Class C amp 1
Q_Q1         2 1 0 Q2
L_L1         2 3  1uH
C_C1         2 3  10nF
R_RL         2 3  60
V_Vdd        3 0 11V
R_Rin        4 1 100
V_Vin        4 0 sin(-1.5 2.7 1591500) DC=-1.5
.model Q2  NPN(Is=14.34f BF=200)

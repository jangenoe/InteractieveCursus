.title opamp
*
* OPAMP MACRO MODEL, SINGLE-POLE 
* connections: non-inverting input
*             | inverting input
*             | |        output
*             | |        |
.subckt opamp 1 2 99 100 6 98
* INPUT IMPEDANCE
RIN 1 2 10MEG
* GAIN BANDWIDTH PRODUCT = 10MHZ
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN 3 0 1 2 100K
RP1 3 4 1K
CP1 4 0 1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER 5 0 4 0 1
ROUT 5 6 10
.ends opamp
* Class C amp 1
Q_Q1         2 1 0 Q2
L_L1         2 3  1uH  
C_C1         2 3  10n  
R_RL         2 3  60  
V_Vdd        3 0 11V
R_Rin        4 1 100
V_Vin        4 5  AC 0.5V 0
V_VinDC      5 0 0.7V
.model Q2  NPN(Is=14.34f BF=200)
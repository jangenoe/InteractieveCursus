.TITLE Transmission Line Example
Rs 1 2 30
O1 2 0 3 0 LOSSYMOD TD=2n
RL 3 0 120
.model LOSSYMOD ltra r=5.14 g=0 l=615E-9 c=246e-12 len=0.0812
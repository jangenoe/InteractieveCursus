Klasse B versterker
*
* SUPPLY VOLTAGES
VPOS 8 0 DC +15V
VNEG 9 0 DC -15V
*
VS2 10 0 DC 0 SIN(0V 5VPEAK 10KHZ)
*
D1  13 10   DNOM
RB1 13 8    10K
Q11 8 13 12 QNPN
*
D2  10 14   DNOM
RB2 14 9    10K
Q12 9 14 12 QPNP
*
RL2 12 0 100
*
* DEVICE MODELS
.model QNPN NPN(BF=50)
.model QPNP PNP(BF=50)
.model DNOM D()

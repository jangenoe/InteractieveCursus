* klasseC   versie2
Q_Q1         2 1 0  Q2
L_L1         0 3    1uH  
C_C1         0 3    10n  
R_R1         0 3    100  
V_V3         4 0    11V
V_V5         1 0    sin(-2 3.09 1591500)
C_C2         2 3    100n  
L_L2         2 4    20uH
.model Q2  NPN(Is=14.34f BF=255.9 Rb=100 )
.title Klasse B versterker  PUSH-PULL PLACED IN OPAMP FEEDBACK LOOP
*
* SUPPLY VOLTAGES
VPOS 8 0 DC +2.5V
VNEG 9 0 DC -2.5V
*
VS3 20 0 DC 0 SIN(0V 1VPEAK 10KHZ)
*
Q21 8 23 22 QNPN
Q22 9 23 22 QPNP
RL3 22 0 100
*
XOpAmp 20 22 8 9 23 8 opamp
*
* DEVICE MODELS
.model QNPN NPN(BF=50)
.model QPNP PNP(BF=50)
.model DNOM D()
Darlington
*
*  PUSH-PULL TRANSISTOR OUTPUT STAGE
Q1 3 1 2 QNPN
Q2 3 2 0 QNPN
*
* DEVICE MODELS
.model QNPN	NPN(BF=50)
* http://www.ecircuitcenter.com/Circuits/smps_buck_vm1/smps_buck_vm1.htm
BUCK_VM1.CIR - BUCK CONVERTER - VOLTAGE MODE CONTROL
* 
* INPUT VOLTAGE
VS	1	0	DC	12
RS	1	2	0.1
*
* BASIC BUCK TOPOLOGY
S1	2 3	11 0 	SW
D1	0	3	DSCH
L1	3	4	50UH
RL1 4	5	0.01
CL	5	6	200UF
R_ESR	6	0	0.1
* MEASURE TOTAL CURRENT OUT W/ RSENSE
RSENSE	5	15	0.01
*
* LOAD
RL	15	0	5
* PULSED LOAD
*ILOAD 15 0	PWL(0US 0A  1000US 0A   1001US 1A  1500US 1A  1501US 0A   2000US 0A)
*
* VOLTAGE MODE CONTROL
* REFERENCE VOLTAGE
VREF	12	0	PWL(0US 0V  10US 0V   201US 5V  1000US 5V)
*
* ERROR AMP AND COMPENSATION
G_ERR	0 10	12 15	0.002
RGAIN	10	0	500K
CGAIN	10	0	10PF
CC	10	7	0.2UF
RC	7	0	2000
DCLAMP	0	10	DZ45
*
* TRIANGLE WAVE FOR PWM 
* (PULSE SOURCE WITH LONG RISE/FALL TIMES)
VTRI	9	0	PULSE(0V 5V 0 4.9US 4.9US 0.1US 10US)
R9	9	0	1MEG
*
* PWM COMPARATOR
ECMP	11	0	TABLE {V(10,9)} = (-5MV 0V) (5MV, 5V) 
R11	11	0	1MEG
*
*
.MODEL	SW	VSWITCH(VON=5V VOFF=0V RON=0.1 ROFF=100K)
.model	DZ45	D( BV=4.5 )
.MODEL DSCH D( IS=0.0002 RS=0.05 CJO=5e-10  )
*
* ANALYSIS
.OPTIONS ABSTOL=1M RELTOL=1M ITL5=0
.TRAN 	1US  	2000US  
*
* VIEW RESULTS
.PRINT	TRAN	V(1) V(15)

.TITLE Transmission Line with driver
MN1 0 1 2 0  NMOS w=150u L=0.50u
MP1 4 1 2 4  PMOS w=350u L=0.50U
VDD 4 0 3.3
O1 2 0 3 0 LOSSYMOD TD=2n
RL 3 0 25
.model LOSSYMOD ltra r=5.14 g=0 l=615E-9 c=246e-12 len=0.1219
.MODEL NMOS NMOS(LEVEL=1 VTO=0.50 KP=90.000E-6 LAMBDA=0.001)
.MODEL PMOS PMOS(LEVEL=1 VTO=-0.45 KP=55.000E-6 LAMBDA=0.001)